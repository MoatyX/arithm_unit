library ieee;
use ieee.std_logic_1164.all;

entity bin_divider is
end bin_divider;
