library ieee;
use ieee.std_logic_1164.all;


entity bin_inverter is
port(
	number: in std_ulogic;
	invertedNumber: out std_ulogic;
);
end bin_inverter;

architecture logic of bin_inverter is
begin
end logic;