library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bin_4bit_divider_test_bench is
end bin_4bit_divider_test_bench;

architecture waveforms of bin_4bit_divider_test_bench is
begin
end waveforms;